﻿{"Id":null,"Data":{"CounterId":"162c2cc0-42cb-4139-a112-ffa6353e1e9a","Timestamp":"2014-05-30T07:18:10.0001613Z","PageSpecificMetrics":null,"Data":0.0,"Id":"8b0b9869-a5d0-46d2-bd0c-04d89b084444"},"Metadata":null}