﻿{"Id":null,"Data":{"CounterId":"0ddeaf92-b1cb-4a32-82cc-b4e0a7f57b01","Timestamp":"2014-05-30T07:20:00.0081594Z","PageSpecificMetrics":{"JsonPageSpecificIntervalHttpLoadStatsByStepUri":{},"JsonPageSpecificLifetimeHttpLoadStatsByStepUri":{},"JsonStatsByStepUri":{}},"Data":null,"Id":"6031bc84-0904-4d0b-b525-acc549d8dbfb"},"Metadata":null}